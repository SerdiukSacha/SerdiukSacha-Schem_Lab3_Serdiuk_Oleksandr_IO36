// ?????????? (?????) ?????? 6-??????? ????????
module ref_sum6bit (
    input  wire [5:0] A,
    input  wire [5:0] B,
    input  wire       cin,
    output wire [5:0] S,
    output wire       cout
);
    assign {cout, S} = A + B + cin;
endmodule

