library verilog;
use verilog.vl_types.all;
entity tb_sum4bit is
end tb_sum4bit;
