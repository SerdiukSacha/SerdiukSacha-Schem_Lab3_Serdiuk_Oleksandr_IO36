library verilog;
use verilog.vl_types.all;
entity tb_sum4bit_basic is
end tb_sum4bit_basic;
