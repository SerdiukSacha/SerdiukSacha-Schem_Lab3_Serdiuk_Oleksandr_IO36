// ?????????? (?????) ?????? 4-??????? ????????
module ref_sum4bit (
    input  wire [3:0] A,
    input  wire [3:0] B,
    input  wire       cin,
    output wire [3:0] S,
    output wire       cout
);
    assign {cout, S} = A + B + cin;
endmodule

