library verilog;
use verilog.vl_types.all;
entity tb_sum6bit is
end tb_sum6bit;
